`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:26:59 11/06/2016 
// Design Name: 
// Module Name:    timer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module select_mode(
    input [3:0] mode,
    input adj_clk_2hz,
    input time_clk_1hz,
    output secondsclk,
    output minutesclk,
    output secondscount,
    output minutescount
    );

    

endmodule
