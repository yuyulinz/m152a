`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:16:42 11/16/2016 
// Design Name: 
// Module Name:    elevtor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module elevtor(
    input [0:7] sw,
    input add,
    input rem,
    input close,
    output [0:3] people,
    output [0:7] floor,
    output dir,
    output open
    );


endmodule
